module vga_record (
    input has_record,
    input [3:0] led1,led2,led3,led4,led5,led6,led7;
    input [9:0] hc,
    input [9:0] vc,
    output has_num
);

parameter hbp        = 144;       //行显示后沿，144（128+16） 96+48
    parameter hfp        = 784;       //行显示前沿784（128+16+640）800-16
    parameter vbp        = 35;       //场显示后延，31（2+29）  ??????? 35(33+2)
    parameter vfp        = 515;     
parameter nums_xs1 = 320;
    parameter nums_xe1 = 340;
    parameter nums_xs2 = 340;
    parameter nums_xe2 = 360;
    parameter nums_xs3 = 360;
    parameter nums_xe3 = 380;
    parameter nums_xs4 = 380;
    parameter nums_xe4 = 400;
    parameter nums_xs5 = 400;
    parameter nums_xe5 = 420;
    parameter nums_xs6 = 420;
    parameter nums_xe6 = 440;
    parameter nums_xs7 = 440;
    parameter nums_xe7 = 460;
    parameter nums_xs8 = 460;
    parameter nums_xe8 = 480;
    parameter nums_ys = 352;
    parameter nums_ye = 416;
    reg [3:0] digit; // stores the digit of current bit
    reg [19:0] words [31:0]; // store the current graph

// 20 x 32
    // 0
parameter [19:0] zero_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00001100000000000000,
    20'b00011100000000000000,
    20'b00111111000000000000,
    20'b01111111000000000000,
    20'b01111111000000000000,
    20'b01110111100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11100001100000000000,
    20'b11100001100000000000,
    20'b11100001100000000000,
    20'b11100001100000000000,
    20'b11100001100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11110011100000000000,
    20'b01110111100000000000,
    20'b01110111100000000000,
    20'b01111111000000000000,
    20'b00111110000000000000
    };
    
    // 1
    parameter [19:0] one_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00001100000000000000,
    20'b00001100000000000000,
    20'b00011100000000000000,
    20'b00111100000000000000,
    20'b00111100000000000000,
    20'b01111100000000000000,
    20'b01111100000000000000,
    20'b01111100000000000000,
    20'b01111100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011110000000000000,
    20'b00011110000000000000,
    20'b00111111000000000000,
    20'b00111111000000000000
    };
    
    // 2
    parameter [19:0] two_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00011100000000000000,
    20'b00011110000000000000,
    20'b00111111000000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b00000011100000000000,
    20'b00000111100000000000,
    20'b00001111100000000000,
    20'b00001111000000000000,
    20'b00001111000000000000,
    20'b00011110000000000000,
    20'b00011110000000000000,
    20'b00111100100000000000,
    20'b00111000100000000000,
    20'b01111001100000000000,
    20'b11111111100000000000,
    20'b11111111100000000000,
    20'b11111111100000000000,
    20'b11111111100000000000
    };
    
    // 3
    parameter [19:0] three_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00001110000000000000,
    20'b00001110000000000000,
    20'b00111111000000000000,
    20'b01111111000000000000,
    20'b01111111000000000000,
    20'b01111111000000000000,
    20'b01100111000000000000,
    20'b01100111000000000000,
    20'b01001111000000000000,
    20'b00001110000000000000,
    20'b00011111100000000000,
    20'b00011111100000000000,
    20'b00011111100000000000,
    20'b00011111100000000000,
    20'b00000011100000000000,
    20'b00000011100000000000,
    20'b00000011100000000000,
    20'b00000011100000000000,
    20'b00000011100000000000,
    20'b11110111100000000000,
    20'b11110111100000000000,
    20'b11111111000000000000,
    20'b11111110000000000000
    };
    
    //4
    parameter [19:0] four_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000011000000000000,
    20'b00000011000000000000,
    20'b00000111000000000000,
    20'b00001111000000000000,
    20'b00001111000000000000,
    20'b00001111000000000000,
    20'b00011111000000000000,
    20'b00011111000000000000,
    20'b00111111000000000000,
    20'b00111111000000000000,
    20'b00111111000000000000,
    20'b01110111000000000000,
    20'b01110111000000000000,
    20'b11110111000000000000,
    20'b11111111110000000000,
    20'b11111111110000000000,
    20'b11111111110000000000,
    20'b11111111110000000000,
    20'b11111111110000000000,
    20'b00000111000000000000,
    20'b00000111000000000000,
    20'b00000111000000000000,
    20'b00000111000000000000
    };
    
    //5
    parameter [19:0] five_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00111111000000000000,
    20'b00111111000000000000,
    20'b00111111000000000000,
    20'b00111111000000000000,
    20'b00111111000000000000,
    20'b00111111000000000000,
    20'b00110000000000000000,
    20'b00110000000000000000,
    20'b00111110000000000000,
    20'b00111110000000000000,
    20'b00111111000000000000,
    20'b00111111100000000000,
    20'b00111111100000000000,
    20'b00111111100000000000,
    20'b00000011100000000000,
    20'b00000011100000000000,
    20'b00000011100000000000,
    20'b00000011100000000000,
    20'b00000011100000000000,
    20'b01110111100000000000,
    20'b01110111100000000000,
    20'b01111111000000000000,
    20'b01111111000000000000
    };
    
    //6
    parameter [19:0] six_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000001000000000000,
    20'b00000011000000000000,
    20'b00001111000000000000,
    20'b00011111000000000000,
    20'b00011111000000000000,
    20'b00111110000000000000,
    20'b00111100000000000000,
    20'b01111100000000000000,
    20'b01111000000000000000,
    20'b01110000000000000000,
    20'b01111111000000000000,
    20'b11111111100000000000,
    20'b11111111100000000000,
    20'b11101111100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11110011100000000000,
    20'b01110111100000000000,
    20'b01110111100000000000,
    20'b01111111100000000000,
    20'b00111111000000000000
    };
    
    //7
    parameter [19:0] seven_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b01111111100000000000,
    20'b11111111100000000000,
    20'b11111111100000000000,
    20'b11111111100000000000,
    20'b11111111100000000000,
    20'b11111111100000000000,
    20'b11000011100000000000,
    20'b11000011100000000000,
    20'b00000111000000000000,
    20'b00000111000000000000,
    20'b00000111000000000000,
    20'b00000110000000000000,
    20'b00000110000000000000,
    20'b00001110000000000000,
    20'b00001110000000000000,
    20'b00001110000000000000,
    20'b00001100000000000000,
    20'b00001100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b00011000000000000000,
    20'b00011000000000000000
    };
    
    //8
    parameter [19:0] eight_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00011110000000000000,
    20'b00011110000000000000,
    20'b00111111000000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b01110011100000000000,
    20'b01110011100000000000,
    20'b01110011100000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b01111111000000000000,
    20'b00111111100000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b01110011100000000000,
    20'b01100001100000000000,
    20'b01110011100000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b00111111000000000000
    };
    
    //9
    parameter [19:0] nine_words[31:0] = {
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00000000000000000000,
    20'b00011100000000000000,
    20'b00011100000000000000,
    20'b01111111000000000000,
    20'b01111111000000000000,
    20'b01111111000000000000,
    20'b11110111100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11100011100000000000,
    20'b11110011100000000000,
    20'b11111111100000000000,
    20'b11111111100000000000,
    20'b01111111100000000000,
    20'b01111111100000000000,
    20'b00111111100000000000,
    20'b00000111100000000000,
    20'b00000111000000000000,
    20'b00001111000000000000,
    20'b00111110000000000000,
    20'b00111110000000000000,
    20'b01111100000000000000,
    20'b01111000000000000000
    };

always @(*) begin
    case (has_record)
        1'b1:
        begin
            if ((hc > = hbp+nums_xs1)&&(hc < hbp+nums_xe1)&&(vc > = vbp+nums_ys)&&(vc < vbp+nums_ye)) begin
                digit = led7;
                has_num = words[vc-vbp-nums_ys][hc-hbp-nums_xs1]
            end else if ((hc > = hbp+nums_xs2)&&(hc < hbp+nums_xe2)&&(vc > = vbp+nums_ys)&&(vc < vbp+nums_ye)) begin
                digit = led6;
                has_num = words[vc-vbp-nums_ys][hc-hbp-nums_xs2]
            end else if ((hc > = hbp+nums_xs3)&&(hc < hbp+nums_xe3)&&(vc > = vbp+nums_ys)&&(vc < vbp+nums_ye)) begin
                digit = led5;
                has_num = words[vc-vbp-nums_ys][hc-hbp-nums_xs3]
            end else if ((hc > = hbp+nums_xs4)&&(hc < hbp+nums_xe4)&&(vc > = vbp+nums_ys)&&(vc < vbp+nums_ye)) begin
                digit = led4;
                has_num = words[vc-vbp-nums_ys][hc-hbp-nums_xs4]
            end else if ((hc > = hbp+nums_xs5)&&(hc < hbp+nums_xe5)&&(vc > = vbp+nums_ys)&&(vc < vbp+nums_ye)) begin
                digit = led3;
                has_num = words[vc-vbp-nums_ys][hc-hbp-nums_xs5]
            end else if ((hc > = hbp+nums_xs6)&&(hc < hbp+nums_xe6)&&(vc > = vbp+nums_ys)&&(vc < vbp+nums_ye)) begin
                digit = led2;
                has_num = words[vc-vbp-nums_ys][hc-hbp-nums_xs6]
            end else if ((hc > = hbp+nums_xs7)&&(hc < hbp+nums_xe7)&&(vc > = vbp+nums_ys)&&(vc < vbp+nums_ye)) begin
                digit = led1;
                has_num = words[vc-vbp-nums_ys][hc-hbp-nums_xs7]
            end else if ((hc > = hbp+nums_xs8)&&(hc < hbp+nums_xe8)&&(vc > = vbp+nums_ys)&&(vc < vbp+nums_ye)) begin
                digit = 0;
                has_num = words[vc-vbp-nums_ys][hc-hbp-nums_xs8]
            end else begin
                has_num=0;
            end
        end 
        default: has_num=0;
    endcase
end    

always @(*) begin
     case (digit)
        4'b0000: words = zero_words;
        4'b0001: words = one_words;
        4'b0010: words = two_words;
        4'b0011: words = three_words;
        4'b0100: words = four_words;
        4'b0101: words = five_words;
        4'b0110: words = six_words;
        4'b0111: words = seven_words;
        4'b1000: words = eight_words;
        4'b1001: words = nine_words;
        default: words = words;
    endcase
end
   
endmodule