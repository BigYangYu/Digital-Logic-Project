//640*480
module vga_top (input clk,
                input debounced_power_on,
                input manul_mode_on,
                input semi_auto_mode_on,
                input auto_mode_on,
                input record,
                input power_now,
                input rst_n,
                output reg hsync,
                output reg vsync,         // hsync and vsync are connected to the port on board.
                   // store the index of horizontal line of current scan position
                output [3:0] red,
                output [3:0] green,
                output [3:0] blue                 // color
                );
     reg [9:0] hc;   // h_cnt
     reg [9:0] vc;  
    reg [3:0] led1,led2,led3,led4,led5,led6,led7;
    reg has_record; // diffe
     reg vsenable; // vertical_sign_enable store the information whether the scan reach an end of a horizontal line
    reg has_word;
    reg has_num; // has word and num store whether the pixel should be lit up.
    wire clk25;
    vga_record record(has_record,led1,led2,led3,led4,led5,led6,led7,hc,vc,has_num) 
    parameter hpixels    = 800;    //行像素点，800
    parameter vlines     = 525;    //行数，521   ???? 525
    parameter hbp        = 144;       //行显示后沿，144（128+16） 96+48
    parameter hfp        = 784;       //行显示前沿784（128+16+640）800-16
    parameter vbp        = 35;       //场显示后延，31（2+29）  ??????? 35(33+2)
    parameter vfp        = 515;       //场显示前沿，511（2+29+480）
    // parameter hpixels = 10'b1100100000;    //行像素点，800
    // parameter vlines  = 10'b1000001101;    //行数，521   ???? 525
    // parameter hbp     = 10'b0010010000;       //行显示后沿，144（128+16） 96+48
    // parameter hfp     = 10'b1100010000;       //行显示前沿784（128+16+640）800-16
    // parameter vbp     = 10'b0000100011;       //场显示后延，31（2+29）  ??????? 35(33+2)
    // parameter vfp     = 10'b0111111111;       //场显示前沿，511（2+29+480）
    parameter cs207_xs   = 160;
    parameter cs207_ys   = 64;
    parameter cs207_xe   = 480;
    parameter cs207_ye   = 128;
    parameter car_xs     = 175;
    parameter car_ys     = 160;
    parameter car_xe     = 465;
    parameter car_ye     = 192;
    parameter name_xs    = 190;
    parameter name_xe    = 450;
    parameter name_ys    = 224;
    parameter name_ye    = 240;
    parameter state_xs   = 160;
    // state_xe depends on the state
    parameter state_ys     = 288;
    parameter state_ye     = 320;
    parameter off_length   = 288;
    parameter manul_length = 352;
    parameter semi_length  = 448;
    parameter auto_length  = 288;
    parameter mileage_xs   = 128;
    parameter mileage_xe   = 320;
    parameter mileage_ys   = 352;
    parameter mileage_ye   = 416;
    parameter nums_xs1 = 320;
    parameter nums_xe1 = 340;
    parameter nums_xs2 = 340;
    parameter nums_xe2 = 360;
    parameter nums_xs3 = 360;
    parameter nums_xe3 = 380;
    parameter nums_xs4 = 380;
    parameter nums_xe4 = 400;
    parameter nums_xs5 = 400;
    parameter nums_xe5 = 420;
    parameter nums_xs6 = 420;
    parameter nums_xe6 = 440;
    parameter nums_xs7 = 440;
    parameter nums_xe7 = 460;
    parameter nums_xs8 = 460;
    parameter nums_xe8 = 480;
    
parameter [0:319] cs207_words[0:63] = {
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000111110000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000111111111111111100000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000011111111111111111111000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000,
    320'b00000000000011111111111111111111111110000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000,
    320'b00000000000111111111111111111111111111000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000,
    320'b00000000001111111111111111111111111111100000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000,
    320'b00000000011111111111111111111111111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000,
    320'b00000000111111111111110000011111111111111000000000000000000000000000011111111111111000011111111111111000000000000000000000000000000011111111111100011111111111100000000000000000000000000000000000000111111111110001111111111100000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000,
    320'b00000001111111111110000000000011111111111000000000000000000000000000011111111110000000000011111111111000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000111111111000000011111111100000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000,
    320'b00000011111111111000000000000000111111111100000000000000000000000000111111111100000000000000111111111100000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000,
    320'b00000011111111110000000000000000011111111100000000000000000000000000111111111000000000000000011111111100000000000000000000000000000111111110000000000000111111111000000000000000000000000000000000001111111100000000000111111110000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000,
    320'b00000111111111100000000000000000001111111110000000000000000000000000111111110000000000000000001111111100000000000000000000000000000111111110000000000000011111111000000000000000000000000000000000001111111100000000000011111111000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000,
    320'b00000111111111000000000000000000001111111110000000000000000000000000111111110000000000000000001111111100000000000000000000000000000111111100000000000000011111111000000000000000000000000000000000011111111000000000000011111111000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000,
    320'b00001111111110000000000000000000000111111111000000000000000000000000111111100000000000000000000111111110000000000000000000000000001111111100000000000000011111111000000000000000000000000000000000011111111000000000000001111111000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000,
    320'b00001111111110000000000000000000000111111111000000000000000000000000111111110000000000000000000111111110000000000000000000000000001111111100000000000000011111111000000000000000000000000000000000011111110000000000000001111111000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000,
    320'b00001111111100000000000000000000000011111100000000000000000000000000111111110000000000000000000111111110000000000000000000000000001111111100000000000000011111111000000000000000000000000000000000011111110000000000000001111111100000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000,
    320'b00011111111100000000000000000000000011000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000111111110000000000000001111111100000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000111111110000000000000001111111100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000111111110000000000000000111111100000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000111111110000000000000000111111100000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000,
    320'b00011111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000,
    320'b00111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000,
    320'b00111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000,
    320'b00111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000,
    320'b00011111110000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000111111100000000000000000111111100000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000,
    320'b00011111111000000000000000000000000001111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000111111110000000000000000111111100000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000,
    320'b00011111111100000000000000000000000011111111000000000000000000000011111111000000000000000000000011111111000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000111111110000000000000001111111100000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000,
    320'b00001111111100000000000000000000000011111111000000000000000000000011111111000000000000000000000011111111000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000111111110000000000000001111111100000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000,
    320'b00001111111100000000000000000000000011111111000000000000000000000011111111000000000000000000000011111111000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000011111110000000000000001111111100000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000,
    320'b00001111111110000000000000000000000111111111000000000000000000000011111111000000000000000000000001111111000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000011111110000000000000001111111000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000,
    320'b00000111111110000000000000000000000111111111000000000000000000000001111111100000000000000000000011111111000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000011111111000000000000001111111000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000,
    320'b00000111111111000000000000000000001111111110000000000000000000000001111111100000000000000000000011111111000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000011111111000000000000011111111000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000,
    320'b00000111111111100000000000000000011111111110000000000000000000000001111111110000000000000000000111111111000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000001111111000000000000011111111000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000,
    320'b00000011111111110000000000000000111111111100000000000000000000000001111111111000000000000000001111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111100000000000111111110000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000,
    320'b00000001111111111000000000000011111111111100000000000000000000000000111111111110000000000000011111111110000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000,
    320'b00000001111111111111000000000111111111111000000000000000000000000000111111111111110000000001111111111100000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000111111111000000011111111100000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000,
    320'b00000000111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000111111111110000111111111100000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000,
    320'b00000000011111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000,
    320'b00000000001111111111111111111111111111000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000,
    320'b00000000000111111111111111111111111110000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000,
    320'b00000000000001111111111111111111111100000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000,
    320'b00000000000000011111111111111111110000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000,
    320'b00000000000000000111111111111110000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    320'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
    };
    
    // a real car
    // 32 x 320 to 290
    parameter [289:0] a_real_car_words[31:0] = {
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000111111110000000000000000000000000000000000000000000111011111000000000000000000000011111100000000000000000000000001111111100000000000000000000111110000000000000000000000000000000000000000000000001111111000000000000000000000000011111111000000000000000000000111011111000000000000000000000,
    290'b00011111111111100000000000000000000000000000000000000001111111111100000000000000000001111111111000000000000000000000111111111111000000000000000000111110000000000000000000000000000000000000000000000011111111110000000000000000000001111111111110000000000000000001111111111100000000000000000000,
    290'b00111111111111110000000000000000000000000000000000000001111111111100000000000000000011111111111100000000000000000001111111111111100000000000000000111110000000000000000000000000000000000000000000001111111111111000000000000000000011111111111111000000000000000001111111111100000000000000000000,
    290'b00111111111111110000000000000000000000000000000000000001111111111000000000000000000111111111111110000000000000000001111111111111100000000000000000111110000000000000000000000000000000000000000000001111111111111100000000000000000011111111111111000000000000000001111111111000000000000000000000,
    290'b01111110000111110000000000000000000000000000000000000001111111111000000000000000001111110000111110000000000000000011111100001111100000000000000000111110000000000000000000000000000000000000000000011111100011111100000000000000000111111000011111000000000000000001111111111000000000000000000000,
    290'b01111100000011110000000000000000000000000000000000000001111110000000000000000000001111100000011111000000000000000011111000000111100000000000000000111110000000000000000000000000000000000000000000011111000001111100000000000000000111110000001111000000000000000001111110000000000000000000000000,
    290'b01111000000011110000000000000000000000000000000000000001111100000000000000000000001111000000011111000000000000000011110000000111100000000000000000111110000000000000000000000000000000000000000000011111000000111100000000000000000111100000001111000000000000000001111100000000000000000000000000,
    290'b00000011111111110000000000000000000000000000000000000001111100000000000000000000001111111111111111000000000000000000000111111111100000000000000000111110000000000000000000000000000000000000000000011110000000000000000000000000000000001111111111000000000000000001111100000000000000000000000000,
    290'b00011111111111110000000000000000000000000000000000000001111100000000000000000000011111111111111111000000000000000000111111111111100000000000000000111110000000000000000000000000000000000000000000011110000000000000000000000000000001111111111111000000000000000001111100000000000000000000000000,
    290'b00111111111111110000000000000000000000000000000000000001111100000000000000000000011111111111111111000000000000000001111111111111100000000000000000111110000000000000000000000000000000000000000000111110000000000000000000000000000011111111111111000000000000000001111100000000000000000000000000,
    290'b01111111111111110000000000000000000000000000000000000001111100000000000000000000011111111111111111000000000000000011111111111111100000000000000000111110000000000000000000000000000000000000000000011110000000000000000000000000000111111111111111000000000000000001111100000000000000000000000000,
    290'b01111110000011110000000000000000000000000000000000000001111100000000000000000000001111000000000000000000000000000011111100000111100000000000000000111110000000000000000000000000000000000000000000011110000000111100000000000000000111111000001111000000000000000001111100000000000000000000000000,
    290'b11111000000011110000000000000000000000000000000000000001111100000000000000000000001111100000011111000000000000000111110000000111100000000000000000111110000000000000000000000000000000000000000000011111000000111100000000000000001111100000001111000000000000000001111100000000000000000000000000,
    290'b11111000000111110000000000000000000000000000000000000001111100000000000000000000001111100000011111000000000000000111110000001111100000000000000000111110000000000000000000000000000000000000000000011111000001111100000000000000001111100000011111000000000000000001111100000000000000000000000000,
    290'b01111100001111110000000000000000000000000000000000000001111100000000000000000000001111111000111111000000000000000011111000011111100000000000000000111110000000000000000000000000000000000000000000011111100011111100000000000000000111110000111111000000000000000001111100000000000000000000000000,
    290'b01111111111111111000000000000000000000000000000000000001111100000000000000000000000111111111111110000000000000000011111111111111110000000000000000111110000000000000000000000000000000000000000000001111111111111000000000000000000111111111111111100000000000000001111100000000000000000000000000,
    290'b01111111111111111000000000000000000000000000000000000001111100000000000000000000000011111111111100000000000000000011111111111111110000000000000000111110000000000000000000000000000000000000000000000111111111111000000000000000000111111111111111100000000000000001111100000000000000000000000000,
    290'b00111111111101111000000000000000000000000000000000000001111100000000000000000000000001111111111000000000000000000001111111111011110000000000000000111110000000000000000000000000000000000000000000000011111111110000000000000000000011111111110111100000000000000001111100000000000000000000000000,
    290'b00001111110000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000111111000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    290'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
    };
    
    0// 260 x 16
    // 12111448 12112323 12112222
    parameter [259:0] sid_words[15:0] = {
    260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    260'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    260'b00110000000111100000001100000000110000000011000000000110000000011000000111000000000000000000110000000111100000001100000000110000000111100000011100000001111000000111000000000000000000110000000111100000001100000000110000000111100000011110000001111000000111100000,
    260'b00110000001111100000001100000000110000000011000000001110000000111000000111100000000000000000110000001111100000001100000000110000001111100000111110000011111000001111100000000000000000110000001111100000001100000000110000001111100000111110000011111000001111100000,
    260'b01110000001111100000011100000001110000000111000000001110000000111000001111100000000000000001110000001111100000011100000001110000001111100000111110000011111000001111100000000000000001110000001111100000011100000001110000001111100000111110000011111000001111100000,
    260'b01110000001101110000011100000001110000000111000000011110000001111000001101100000000000000001110000001101110000011100000001110000001101110000110110000011011100001101100000000000000001110000001101110000011100000001110000001101110000110111000011011100001101110000,
    260'b01110000001101110000011100000001110000000111000000011110000001111000001111100000000000000001110000001101110000011100000001110000001101110000110110000011011100001101100000000000000001110000001101110000011100000001110000001101110000110111000011011100001101110000,
    260'b01110000000001100000011100000001110000000111000000011110000001111000001111100000000000000001110000000001100000011100000001110000000001100000001110000000011000000011100000000000000001110000000001100000011100000001110000000001100000000110000000011000000001100000,
    260'b00110000000011100000001100000000110000000011000000111110000011111000001111100000000000000000110000000011100000001100000000110000000011100000001110000000111000000011100000000000000000110000000011100000001100000000110000000011100000001110000000111000000011100000,
    260'b00110000000111100000001100000000110000000011000000111111000011111100001111110000000000000000110000000111100000001100000000110000000111100000001111000001111000000011110000000000000000110000000111100000001100000000110000000111100000011110000001111000000111100000,
    260'b00110000000111000000001100000000110000000011000000111111000011111100001101110000000000000000110000000111000000001100000000110000000111000000110111000001110000001101110000000000000000110000000111000000001100000000110000000111000000011100000001110000000111000000,
    260'b00110000001111000000001100000000110000000011000000111111000011111100001100110000000000000000110000001111000000001100000000110000001111000000110111000011110000001101110000000000000000110000001111000000001100000000110000001111000000111100000011110000001111000000,
    260'b00110000001111110000001100000000110000000011000000000110000000011000001111110000000000000000110000001111110000001100000000110000001111110000111111000011111100001111110000000000000000110000001111110000001100000000110000001111110000111111000011111100001111110000,
    260'b00110000001111110000001100000000110000000011000000000110000000011000001111100000000000000000110000001111110000001100000000110000001111110000111110000011111100001111100000000000000000110000001111110000001100000000110000001111110000111111000011111100001111110000,
    260'b00110000001111110000001100000000110000000011000000000110000000011000000111100000000000000000110000001111110000001100000000110000001111110000011110000011111100000111100000000000000000110000001111110000001100000000110000001111110000111111000011111100001111110000,
    260'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
    };
    
    // power off
    // 288 x 32
    parameter [287:0] power_off_words[31:0] = {
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000001111111000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000011111111000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000111111111000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000111110000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b001110011111100000000000000000000000011111110000000000000000000011110000011111000001111000000000000000111111000000000000000000000011101111100000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111110000000000000000000000011111111100000000000000000000000,
    288'b011111111111110000000000000000000000111111111100000000000000000111110000011111000001111100000000000011111111110000000000000000000111111111110000000000000000000000000000000000000000000000000000000011111111110000000000000000001111111111000000000000000000000011111111110000000000000000000000,
    288'b011111111111111000000000000000000011111111111110000000000000000011110000011111000001111000000000000111111111111000000000000000000111111111110000000000000000000000000000000000000000000000000000001111111111111000000000000000001111111111000000000000000000000011111111110000000000000000000000,
    288'b011111111111111100000000000000000011111111111111000000000000000011111000011111100011111000000000001111111111111100000000000000000111111111100000000000000000000000000000000000000000000000000000001111111111111100000000000000001111111111000000000000000000000011111111110000000000000000000000,
    288'b011111110001111100000000000000000111111000111111100000000000000011111000111111100011111000000000011111100001111100000000000000000111111111100000000000000000000000000000000000000000000000000000011111100011111110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111100000111110000000000000000111110000001111100000000000000011111000111111100011110000000000011111000000111110000000000000000111111000000000000000000000000000000000000000000000000000000000011111000000111110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111000000111110000000000000000111100000001111100000000000000001111000111111100011110000000000011110000000111110000000000000000111110000000000000000000000000000000000000000000000000000000000011110000000111110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111000000011110000000000000001111100000000111100000000000000001111101111111110111110000000000011111111111111110000000000000000111110000000000000000000000000000000000000000000000000000000000111110000000011110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111000000011110000000000000001111100000000111100000000000000001111101111111110111110000000000111111111111111110000000000000000111110000000000000000000000000000000000000000000000000000000000111110000000011110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011110000000011110000000000000001111100000000111100000000000000000111101111011110111100000000000111111111111111110000000000000000111110000000000000000000000000000000000000000000000000000000000111110000000011110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111000000011110000000000000001111100000000111100000000000000000111111111011111111100000000000111111111111111110000000000000000111110000000000000000000000000000000000000000000000000000000000111110000000011110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111000000011110000000000000000111100000000111100000000000000000111111111011111111100000000000011110000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000011110000000011110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111000000111110000000000000000111110000001111100000000000000000011111110011111111000000000000011111000000111110000000000000000111110000000000000000000000000000000000000000000000000000000000011111000000111110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111100000111110000000000000000111110000001111100000000000000000011111110001111111000000000000011111000000111110000000000000000111110000000000000000000000000000000000000000000000000000000000011111000000111110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111110011111100000000000000000111111000111111100000000000000000011111110001111111000000000000011111110001111110000000000000000111110000000000000000000000000000000000000000000000000000000000011111100011111110000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111111111111100000000000000000011111111111111000000000000000000001111110001111110000000000000001111111111111100000000000000000111110000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111111111111000000000000000000011111111111110000000000000000000001111100001111110000000000000000111111111111000000000000000000111110000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111111111110000000000000000000000111111111100000000000000000000001111100000111110000000000000000011111111110000000000000000000111110000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011110000000000000000000000000000111100000000000000000000000000,
    288'b011111011111000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
    };
    
    
    // manul mode
    // 352x32
    parameter [351:0] manul_mode_words[31:0] = {
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    352'b0011100111110000011111100000000000000111111110000000000000000000001110011111100000000000000000000011100000001111000000000000000000000111111110000000000000000000011111000000000000000000000000000000000000000000000000000000000000111001111100000111111000000000000001111111000000000000000000000000011111101111000000000000000000000011111100000000000000000000,
    352'b0111111111111101111111110000000000011111111111100000000000000000011111111111111000000000000000000111110000001111000000000000000000011111111111100000000000000000011111000000000000000000000000000000000000000000000000000000000001111111111111011111111100000000000011111111110000000000000000000001111111111111000000000000000000001111111111000000000000000000,
    352'b0111111111111111111111111000000000111111111111110000000000000000011111111111111100000000000000000111110000001111000000000000000000111111111111110000000000000000011111000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000001111111111111000000000000000000011111111111111000000000000000000011111111111100000000000000000,
    352'b0111111111111111111111111000000000111111111111110000000000000000011111111111111100000000000000000111110000001111000000000000000000111111111111110000000000000000011111000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000001111111111111100000000000000000011111111111111000000000000000000111111111111110000000000000000,
    352'b0111111100111111110011111000000001111110000111110000000000000000011111110001111100000000000000000111110000001111000000000000000001111110000111110000000000000000011111000000000000000000000000000000000000000000000000000000000001111111001111111100111110000000011111100011111110000000000000000111111000111111000000000000000001111110000111110000000000000000,
    352'b0111111000011111000001111000000001111100000011110000000000000000011111100001111100000000000000000111110000001111000000000000000001111100000011110000000000000000011111000000000000000000000000000000000000000000000000000000000001111110000111110000011110000000011111000000111110000000000000000111110000011111000000000000000001111100000011111000000000000000,
    352'b0111110000011111000001111000000001111000000011110000000000000000011111000000111100000000000000000111110000001111000000000000000001111000000011110000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000011110000000111110000000000000000111100000011111000000000000000001111000000011111000000000000000,
    352'b0111110000011111000001111000000000000011111111110000000000000000011111000000111100000000000000000111110000001111000000000000000000000011111111110000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000001111111111111111000000000000000,
    352'b0111110000011111000001111000000000011111111111110000000000000000011111000000111100000000000000000111110000001111000000000000000000011111111111110000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000011111111111111111000000000000000,
    352'b0111110000011111000001111000000000111111111111110000000000000000011111000000111100000000000000000111110000001111000000000000000000111111111111110000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000011111111111111111000000000000000,
    352'b0111110000011111000001111000000001111111111111110000000000000000011111000000111100000000000000000111110000001111000000000000000001111111111111110000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000011111111111111111000000000000000,
    352'b0111110000011111000001111000000001111110000011110000000000000000011111000000111100000000000000000111110000001111000000000000000001111110000011110000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000011110000000011110000000000000001111100000001111000000000000000001111000000000000000000000000000,
    352'b0111110000011111000001111000000011111000000011110000000000000000011111000000111100000000000000000111110000001111000000000000000011111000000011110000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000011111000000111110000000000000000111110000011111000000000000000001111100000011111000000000000000,
    352'b0111110000011111000001111000000011111000000111110000000000000000011111000000111100000000000000000111110000011111000000000000000011111000000111110000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000011111000000111110000000000000000111110000011111000000000000000001111100000011111000000000000000,
    352'b0111110000011111000001111000000001111100001111110000000000000000011111000000111100000000000000000111111001111111000000000000000001111100001111110000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000011111100011111110000000000000000111111000111111000000000000000001111111000111111000000000000000,
    352'b0111110000011111000001111000000001111111111111111000000000000000011111000000111100000000000000000011111111111111000000000000000001111111111111111000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000001111111111111100000000000000000011111111111111000000000000000000111111111111110000000000000000,
    352'b0111110000011111000001111000000001111111111111111000000000000000011111000000111100000000000000000011111111111111000000000000000001111111111111111000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000001111111111111000000000000000000011111111111111000000000000000000011111111111100000000000000000,
    352'b0111110000011111000001111000000000111111111101111000000000000000011111000000111100000000000000000001111111111111000000000000000000111111111101111000000000000000011111000000000000000000000000000000000000000000000000000000000001111100000111110000011110000000000011111111110000000000000000000000111111111111000000000000000000001111111111000000000000000000,
    352'b0000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000011111000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000011111000000000000000000000000000011111100000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    352'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
    };
    
    
    // semi-auto mode
    // 448x32
    parameter [447:0] semi_auto_mode_words[31:0] = {
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    448'b0000111111100000000000000000000000000011111100000000000000000000001110011111000001111110000000000011100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000011100000001111000000000000000011111111100000000000000000000000000001111111000000000000000000000000000000000000000000000000000000111001111100000111111000000000000001111111000000000000000000000000011111101111000000000000000000000011111100000000000000000000,
    448'b0011111111111000000000000000000000001111111111000000000000000000011111111111110111111111000000000111110000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000111110000001111000000000000000011111111100000000000000000000000000011111111110000000000000000000000000000000000000000000000000001111111111111011111111100000000000011111111110000000000000000000001111111111111000000000000000000001111111111000000000000000000,
    448'b0111111111111100000000000000000000011111111111100000000000000000011111111111111111111111100000000111110000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000111110000001111000000000000000011111111100000000000000000000000001111111111111000000000000000000000000000000000000000000000000001111111111111111111111110000000001111111111111000000000000000000011111111111111000000000000000000011111111111100000000000000000,
    448'b0111111111111100000000000000000000111111111111110000000000000000011111111111111111111111100000000111110000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000111110000001111000000000000000011111111100000000000000000000000001111111111111100000000000000000000000000000000000000000000000001111111111111111111111110000000001111111111111100000000000000000011111111111111000000000000000000111111111111110000000000000000,
    448'b0111110001111110000000000000000001111110000111110000000000000000011111110011111111001111100000000111110000000000000000000000000000000000000000000000000000000000011111100001111100000000000000000111110000001111000000000000000000111100000000000000000000000000011111100011111110000000000000000000000000000000000000000000000001111111001111111100111110000000011111100011111110000000000000000111111000111111000000000000000001111110000111110000000000000000,
    448'b0111100000111110000000000000000001111100000011111000000000000000011111100001111100000111100000000111110000000000000000000000000000000000000000000000000000000000011111000000111100000000000000000111110000001111000000000000000000111100000000000000000000000000011111000000111110000000000000000000000000000000000000000000000001111110000111110000011110000000011111000000111110000000000000000111110000011111000000000000000001111100000011111000000000000000,
    448'b0111111000010000000000000000000001111000000011111000000000000000011111000001111100000111100000000111110000000000000000000000000000000000000000000000000000000000011110000000111100000000000000000111110000001111000000000000000000111100000000000000000000000000011110000000111110000000000000000000000000000000000000000000000001111100000111110000011110000000011110000000111110000000000000000111100000011111000000000000000001111000000011111000000000000000,
    448'b0111111111100000000000000000000001111111111111111000000000000000011111000001111100000111100000000111110000000000000000000000000011111111110000000000000000000000000000111111111100000000000000000111110000001111000000000000000000111100000000000000000000000000111110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000001111111111111111000000000000000,
    448'b0111111111111000000000000000000011111111111111111000000000000000011111000001111100000111100000000111110000000000000000000000000011111111110000000000000000000000000111111111111100000000000000000111110000001111000000000000000000111100000000000000000000000000111110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000011111111111111111000000000000000,
    448'b0011111111111110000000000000000011111111111111111000000000000000011111000001111100000111100000000111110000000000000000000000000011111111110000000000000000000000001111111111111100000000000000000111110000001111000000000000000000111100000000000000000000000000111110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000011111111111111111000000000000000,
    448'b0000111111111110000000000000000011111111111111111000000000000000011111000001111100000111100000000111110000000000000000000000000011111111110000000000000000000000011111111111111100000000000000000111110000001111000000000000000000111100000000000000000000000000111110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000011111111111111111000000000000000,
    448'b0000000011111110000000000000000001111000000000000000000000000000011111000001111100000111100000000111110000000000000000000000000011111111110000000000000000000000011111100000111100000000000000000111110000001111000000000000000000111100000000000000000000000000011110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000011110000000011110000000000000001111100000001111000000000000000001111000000000000000000000000000,
    448'b1111100000111111000000000000000001111100000011111000000000000000011111000001111100000111100000000111110000000000000000000000000000000000000000000000000000000000111110000000111100000000000000000111110000001111000000000000000000111100000000000000000000000000011111000000111110000000000000000000000000000000000000000000000001111100000111110000011110000000011111000000111110000000000000000111110000011111000000000000000001111100000011111000000000000000,
    448'b1111100000011111000000000000000001111100000011111000000000000000011111000001111100000111100000000111110000000000000000000000000000000000000000000000000000000000111110000001111100000000000000000111110000011111000000000000000000111100000000000000000000000000011111000000111110000000000000000000000000000000000000000000000001111100000111110000011110000000011111000000111110000000000000000111110000011111000000000000000001111100000011111000000000000000,
    448'b0111110000111110000000000000000001111111000111111000000000000000011111000001111100000111100000000111110000000000000000000000000000000000000000000000000000000000011111000011111100000000000000000111111001111111000000000000000000111111000000000000000000000000011111100011111110000000000000000000000000000000000000000000000001111100000111110000011110000000011111100011111110000000000000000111111000111111000000000000000001111111000111111000000000000000,
    448'b0111111111111110000000000000000000111111111111110000000000000000011111000001111100000111100000000111110000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000011111111111111000000000000000000111111100000000000000000000000001111111111111100000000000000000000000000000000000000000000000001111100000111110000011110000000001111111111111100000000000000000011111111111111000000000000000000111111111111110000000000000000,
    448'b0011111111111100000000000000000000011111111111100000000000000000011111000001111100000111100000000111110000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000011111111111111000000000000000000111111100000000000000000000000001111111111111000000000000000000000000000000000000000000000000001111100000111110000011110000000001111111111111000000000000000000011111111111111000000000000000000011111111111100000000000000000,
    448'b0011111111111000000000000000000000001111111111000000000000000000011111000001111100000111100000000111110000000000000000000000000000000000000000000000000000000000001111111111011110000000000000000001111111111111000000000000000000011111100000000000000000000000000011111111110000000000000000000000000000000000000000000000000001111100000111110000011110000000000011111111110000000000000000000000111111111111000000000000000000001111111111000000000000000000,
    448'b0000011111100000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000011111000000000000000000000000001111100000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000011111000000000000000000000000000011111100000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
    };
    
    
    // auto mode
    // 288x32
    parameter [287:0] auto_mode_words[31:0] = {
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000,
    288'b000001111111100000000000000000000011100000001111000000000000000011111111100000000000000000000000000001111111000000000000000000000000000000000000000000000000000000111001111100000111111000000000000001111111000000000000000000000000011111101111000000000000000000000011111100000000000000000000,
    288'b000111111111111000000000000000000111110000001111000000000000000011111111100000000000000000000000000011111111110000000000000000000000000000000000000000000000000001111111111111011111111100000000000011111111110000000000000000000001111111111111000000000000000000001111111111000000000000000000,
    288'b001111111111111100000000000000000111110000001111000000000000000011111111100000000000000000000000001111111111111000000000000000000000000000000000000000000000000001111111111111111111111110000000001111111111111000000000000000000011111111111111000000000000000000011111111111100000000000000000,
    288'b001111111111111100000000000000000111110000001111000000000000000011111111100000000000000000000000001111111111111100000000000000000000000000000000000000000000000001111111111111111111111110000000001111111111111100000000000000000011111111111111000000000000000000111111111111110000000000000000,
    288'b011111100001111100000000000000000111110000001111000000000000000000111100000000000000000000000000011111100011111110000000000000000000000000000000000000000000000001111111001111111100111110000000011111100011111110000000000000000111111000111111000000000000000001111110000111110000000000000000,
    288'b011111000000111100000000000000000111110000001111000000000000000000111100000000000000000000000000011111000000111110000000000000000000000000000000000000000000000001111110000111110000011110000000011111000000111110000000000000000111110000011111000000000000000001111100000011111000000000000000,
    288'b011110000000111100000000000000000111110000001111000000000000000000111100000000000000000000000000011110000000111110000000000000000000000000000000000000000000000001111100000111110000011110000000011110000000111110000000000000000111100000011111000000000000000001111000000011111000000000000000,
    288'b000000111111111100000000000000000111110000001111000000000000000000111100000000000000000000000000111110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000001111111111111111000000000000000,
    288'b000111111111111100000000000000000111110000001111000000000000000000111100000000000000000000000000111110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000011111111111111111000000000000000,
    288'b001111111111111100000000000000000111110000001111000000000000000000111100000000000000000000000000111110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000011111111111111111000000000000000,
    288'b011111111111111100000000000000000111110000001111000000000000000000111100000000000000000000000000111110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000111110000000011110000000000000001111100000001111000000000000000011111111111111111000000000000000,
    288'b011111100000111100000000000000000111110000001111000000000000000000111100000000000000000000000000011110000000011110000000000000000000000000000000000000000000000001111100000111110000011110000000011110000000011110000000000000001111100000001111000000000000000001111000000000000000000000000000,
    288'b111110000000111100000000000000000111110000001111000000000000000000111100000000000000000000000000011111000000111110000000000000000000000000000000000000000000000001111100000111110000011110000000011111000000111110000000000000000111110000011111000000000000000001111100000011111000000000000000,
    288'b111110000001111100000000000000000111110000011111000000000000000000111100000000000000000000000000011111000000111110000000000000000000000000000000000000000000000001111100000111110000011110000000011111000000111110000000000000000111110000011111000000000000000001111100000011111000000000000000,
    288'b011111000011111100000000000000000111111001111111000000000000000000111111000000000000000000000000011111100011111110000000000000000000000000000000000000000000000001111100000111110000011110000000011111100011111110000000000000000111111000111111000000000000000001111111000111111000000000000000,
    288'b011111111111111110000000000000000011111111111111000000000000000000111111100000000000000000000000001111111111111100000000000000000000000000000000000000000000000001111100000111110000011110000000001111111111111100000000000000000011111111111111000000000000000000111111111111110000000000000000,
    288'b011111111111111110000000000000000011111111111111000000000000000000111111100000000000000000000000001111111111111000000000000000000000000000000000000000000000000001111100000111110000011110000000001111111111111000000000000000000011111111111111000000000000000000011111111111100000000000000000,
    288'b001111111111011110000000000000000001111111111111000000000000000000011111100000000000000000000000000011111111110000000000000000000000000000000000000000000000000001111100000111110000011110000000000011111111110000000000000000000000111111111111000000000000000000001111111111000000000000000000,
    288'b000011111100000000000000000000000000011111000000000000000000000000001111100000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000011111000000000000000000000000000011111100000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    288'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
    };
    
    
    // mileage
    // 199 x 32  from 224
    // 192 = 32*6
    parameter [191:0] mileage_words[31:0] = {
    192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000111110000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000111110000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000111110000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000111110000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000111110000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
    192'b001110011111000001111110000000000011100000000000000111110000000000000000000111111000000000000000000000001111111100000000000000000000001111110011100000000000000000000011111100000000000000000000,
    192'b011111111111110111111111000000000111110000000000000111110000000000000000011111111110000000000000000000111111111111000000000000000000111111111111100000000000000000001111111111000000000000000000,
    192'b011111111111111111111111100000000111110000000000000111110000000000000000111111111111000000000000000001111111111111100000000000000001111111111111100000000000000000011111111111100000000000000000,
    192'b011111111111111111111111100000000111110000000000000111110000000000000001111111111111100000000000000001111111111111100000000000000001111111111111100000000000000000111111111111110000000000000000,
    192'b011111110011111111001111100000000111110000000000000111110000000000000011111100001111100000000000000011111100001111100000000000000011111100011111100000000000000001111110000111110000000000000000,
    192'b011111100001111100000111100000000111110000000000000111110000000000000011111000000111110000000000000011111000000111100000000000000011111000001111100000000000000001111100000011111000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000011110000000111110000000000000011110000000111100000000000000111110000000111100000000000000001111000000011111000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000011111111111111110000000000000000000111111111100000000000000111110000000111100000000000000001111111111111111000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000111111111111111110000000000000000111111111111100000000000000111110000000111100000000000000011111111111111111000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000111111111111111110000000000000001111111111111100000000000000111110000000111100000000000000011111111111111111000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000111111111111111110000000000000011111111111111100000000000000111110000000111100000000000000011111111111111111000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000011110000000000000000000000000011111100000111100000000000000011110000000111100000000000000001111000000000000000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000011111000000111110000000000000111110000000111100000000000000011111000001111100000000000000001111100000011111000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000011111000000111110000000000000111110000001111100000000000000011111000001111100000000000000001111100000011111000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000011111110001111110000000000000011111000011111100000000000000011111110111111100000000000000001111111000111111000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000001111111111111100000000000000011111111111111110000000000000001111111111111100000000000000000111111111111110000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000000111111111111000000000000000011111111111111110000000000000000111111111111100000000000000000011111111111100000000000000000,
    192'b011111000001111100000111100000000111110000000000000111110000000000000000011111111110000000000000000001111111111011110000000000000000011111111111100000000000000000001111111111000000000000000000,
    192'b000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000011111100000000000000000000011000000000111100000000000000000000011111100000000000000000000,
    192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001111100000000000000000000000000000000000000000000000,
    192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000001111100000000000000000000000000000000000000000000000
    };
    
   
    always@(posedge clk)
    begin
        clk25 <= ~clk25;
    end
    
    always @(posedge clk25) begin
        if (hc == hpixels - 1)
        begin
            hc       <= 0;
            vsenable <= 1;
        end
        else
        begin
            hc       <= hc +1;
            vsenable <= 0;
        end
    end
    
    always @(*) begin
        if (hc < 96)  //同步为96 96 is the sync time
            hsync = 0;
        else
            hsync = 1;
    end
    
    // update the index of current vertical line when the scan reach the end of a horizontal line
    always @(posedge clk25) begin
        if (vsenable == 1) // when the scan reach the end of a horizontal line
        begin
            if (vc == vlines - 1)
                vc <= 0;
            else
                vc <= vc + 1;
        end
        else
            vc <= vc;
    end
    
    
    always @(*) begin
        if (vc < 2)   //同步为2  2 is the sync time
            vsync = 0;
        else
            vsync = 1;
    end
    
   
    
    //     (hc > = hbp+)&&(hc < hbp+)&&(vc > = vbp+)&&(vc < vbp+)
    // always @(*) begin
    //     if (((hc > = hbp+cs207_xs)&&(hc < hbp+cs207_xe)&&(vc > = vbp+cs207_ys)&&(vc < vbp+cs207_ye))||
    //     ((hc > = hbp+car_xs)&&(hc < hbp+car_xe)&&(vc > = vbp+car_ys)&&(vc < vbp+car_ye))||
    //     ((hc > = hbp+name_xs)&&(hc < hbp+name_xe)&&(vc > = vbp+name_ys)&&(vc < vbp+name_ye)))
    //     begin
    //         has_word = 1'b1;
    //     end
    //     else
    //     begin
    //        casex (debounced_power_on)
    //         0: // power_off
    //         begin
    //             if ((hc > = hbp+state_xs)&&(hc < hbp+state_xs+off_length)&&(vc > = vbp+state_ys)&&(vc < vbp+state_ye))
    //         end
    //         default:
    //     endcase
    //     end
    // end
    
    always @(*) begin
        casex (debounced_power_on)
            0: begin
                if ((hc > = hbp+state_xs)&&(hc < hbp+state_xs+off_length)&&(vc > = vbp+state_ys)&&(vc < vbp+state_ye))
                begin
                    has_word = power_off_words[vc-vbp-state_ys][hc-hbp-state_xs:hc-hbp-state_xs];
                end
                else
                begin
                    has_word = 0;
                end
            end
            default: begin
                case ({manul_mode_on,semi_auto_mode_on,auto_mode_on})
                    3'b100:
                    begin
                        if ((hc > = hbp+state_xs)&&(hc < hbp+state_xs+manul_length)&&(vc > = vbp+state_ys)&&(vc < vbp+state_ye))
                        begin
                            has_word = power_off_words[vc-vbp-state_ys][hc-hbp-state_xs:hc-hbp-state_xs];
                            has_record =0;
                        end
                        else
                        begin
                            if (rst_n&&power_now) begin
                                // led7 = 0; //0
                                // led6 = 0; //0
                                // led5 = 0; //0
                                // led4 = 0; //0
                                // led3 = 0; //0
                                // led2 = 0; //0
                                // led1 = 0; //0
                                has_word=0;
                                has_record = 0;
                            end
                            else begin
                                led7 = (record/100_0000)%10;
                                led6 = (record/10_0000)%10;
                                led5 = (record/1_0000)%10;
                                led4 = (record/1_000)%10;
                                led3 = (record/100)%10;
                                led2 = (record/10)%10;
                                led1 = record%10;
                                has_word=0;
                                has_record =1;
                            end
                        end
                    end
                    3'b010:
                    begin
                        has_record = 0;
                        if ((hc > = hbp+state_xs)&&(hc < hbp+state_xs+semi_length)&&(vc > = vbp+state_ys)&&(vc < vbp+state_ye))
                        begin
                            has_word = power_off_words[vc-vbp-state_ys][hc-hbp-state_xs:hc-hbp-state_xs];
                        end
                        else
                        begin
                            has_word = 0;
                        end
                    end
                    3'b001:
                    begin
                        has_record = 0;
                        if ((hc > = hbp+state_xs)&&(hc < hbp+state_xs+auto_length)&&(vc > = vbp+state_ys)&&(vc < vbp+state_ye))
                        begin
                            has_word = power_off_words[vc-vbp-state_ys][hc-hbp-state_xs:hc-hbp-state_xs];
                        end
                        else
                        begin
                            has_word = 0;
                        end
                    end
                    default:begin
                        has_word = 0;
                        has_word = 0;
                    end 
                endcase
            end
        endcase
    end
    
    always @(*) begin // this block control color
        red   = 0;   //这里三个置零起到消隐作用
        blue  = 0;
        green = 0;
        case ({has_word,has_num})
            1'b1:
            begin   //白色
                red   = 4'b1111;
                green = 4'b1111;
                blue  = 4'b1111;
            end
            default:
            begin
                red   = 0;   //这里三个置零起到消隐作用
                blue  = 0;
                green = 0;
            end
        endcase
    end
endmodule
    
    
    
    
    
    
    
